b0VIM 7.2      H�nLP�8_D  foca                                    dalek.local                             ~foca/Projects/cubox/datacatalog-web/app/models                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              utf-8	U3210    #"! U                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 tp                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        ad  Y  �            �  c  )    �  [      �  �  �  �  �  �  �  l  _  L  ;  #                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                006ÿuser_session.rb 006ÿu006ÿuser_session.rb 006006ÿuser_session006ÿuser_session.r006ÿuser_ses006ÿuser_session.rb 006ÿuser006ÿ006ÿ006ÿ006ÿ006ÿ006ÿ006ÿuser_session.rb user.rb submission.rb notifier.rb data_suggestion.rb contact_submission.rb ../ " ============================================================================ "   Quick Help: <F1>:help  -:go up dir  D:delete  R:rename  s:sort-by  x:exec "   Sort sequence: [\/]$,\<core\%(\.\d\+\)\=\>,\.h$,\.c$,\.cpp$,*,\.o$,\.obj$,\.info$,\.swp$,\.bak$,\~$ "   Sorted by      name "   /Users/foca/Projects/cubox/datacatalog-web/app/models " Netrw Directory Listing                                        (netrw v136) " ============================================================================ 